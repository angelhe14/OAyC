library ieee;
use ieee.std_logic_1164.all;

entity register3x is 
	port( CLK: in std_logic;
				RESET: in std_logic;
			ENTRADA: in std_logic_vector(2 downto 0);
			SALIDA: out std_logic_vector(2 downto 0));
end register3X;

architecture behavioral of register3x is
signal internal_value: std_logic_vector (2 downto 0):= B"000";
begin
	process (CLK, RESET, ENTRADA)
	begin
		if RESET = '0' then
			internal_value <= B"000";
		elsif rising_edge (CLK) then
			internal_value <= ENTRADA;
		end if;
	end process;
	
	process (internal_value)
	begin
		SALIDA<= internal_value;
	end process;
end behavioral;